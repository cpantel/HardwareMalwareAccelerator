`timescale 1ns/1ps

module uart_testbench;
  reg simul_Clock;
  reg send;
  wire active;
  wire done;
  wire tx;

localparam char = 8'b10100011;

  initial begin
    simul_Clock = 1'b0;
    forever simul_Clock = #2.5 ~simul_Clock;
  end

  initial begin
    send = 1'b0;
    #100 send = 1'b1;
    #10 send = 1'b0;
    
  end

  initial begin
    repeat(64) @(negedge simul_Clock);
    $finish;
  end

uart_tx uart_tx(
   .i_Clock(simul_Clock),
   .i_Tx_DV(send),
   .i_Tx_Byte(char),
   .o_Tx_Active(active),
   .o_Tx_Serial(tx),
   .o_Tx_Done(done)
);

endmodule
